`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Create Date:    Tue May 07 14:31:56 2013
// Design Name: 
// Module Name:    netlist_1_EMPTY
//////////////////////////////////////////////////////////////////////////////////
module netlist_1_EMPTY(sensor, servo, seg, led, an, clk, reset, rx, tx);
  input [2:0] sensor;
  output [1:0] servo;
  output [7:0] seg;
  output [7:0] led;
  output [3:0] an;
  input clk;
  input reset;
  input rx;
  output tx;


endmodule
